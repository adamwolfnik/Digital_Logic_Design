module AND_gate(a,b,y);
input a,b;
output y;
and A1(y,a,b);
endmodule;

